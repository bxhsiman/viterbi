//==============================================================================
// 文件名: viterbi_encode9.v
// 描述: Viterbi编码器模块 (Viterbi Encoder)
//
// 模块功能和原理:
// 1. 实现(2,1,8)卷积编码器，约束长度为9
// 2. 使用两个生成多项式产生两路编码输出
// 3. 编码率为1/2，即每个输入位产生2个输出位
//
// 编码参数:
// - 约束长度K=9 (需要8个存储单元)
// - 编码率R=1/2 (1位输入，2位输出)
// - 生成多项式:
//   * G1 = 110101111 (八进制557)
//   * G2 = 100011101 (八进制435)
//
// 工作原理:
// 1. 输入数据X通过8级移位寄存器(ShReg)
// 2. 两个生成多项式分别与移位寄存器内容进行按位与运算
// 3. 对与运算结果进行异或运算，得到编码输出
// 4. 输出经过D触发器同步后输出Y[1:0]
//
// 数据流:
// X → ShReg[8:0] → PolyA&ShReg / PolyB&ShReg → XOR → Y[1:0]
//==============================================================================

//==============================================================================
// 模块名: viterbi_encode9
// 功能: (2,1,8)卷积编码器，实现1/2编码率的卷积编码
// 输入:
//   - X: 输入数据位
//   - Clock: 时钟信号
//   - Reset: 复位信号
// 输出:
//   - Y: 2位编码输出[Y1, Y0]
//==============================================================================
module viterbi_encode9(X,Y,Clock,Reset); 

// 端口定义
input X, Clock, Reset;                        // 输入信号
output [1:0] Y;                               // 编码输出

// 内部信号定义
wire [1:0] Yt;                                // 编码结果(未同步)
wire X, Clock, Reset;                         // 输入信号重声明

wire [8:0] PolyA, PolyB;                      // 生成多项式
wire [8:0] wA, wB, ShReg;                     // 中间计算信号

   //===========================================================================
   // 生成多项式定义
   // G1 = 110101111 (八进制557) - 对应Y[1]输出
   // G2 = 100011101 (八进制435) - 对应Y[0]输出
   //===========================================================================
   assign   PolyA = 9'b110_101_111;           // 生成多项式A (G1)
   assign   PolyB = 9'b100_011_101;           // 生成多项式B (G2)

   //===========================================================================
   // 卷积运算
   // 将移位寄存器内容与生成多项式进行按位与运算
   //===========================================================================
   assign wA = PolyA & ShReg;                 // 多项式A的卷积结果
   assign wB = PolyB & ShReg;                 // 多项式B的卷积结果

   //===========================================================================
   // 8级移位寄存器实现
   // ShReg[8]为当前输入，ShReg[7:0]为历史数据
   //===========================================================================
   assign ShReg[8] = X;                       // 当前输入位
   pDFF dff7(ShReg[8], ShReg[7], Clock, Reset); // 第7级D触发器
   pDFF dff6(ShReg[7], ShReg[6], Clock, Reset); // 第6级D触发器  
   pDFF dff5(ShReg[6], ShReg[5], Clock, Reset); // 第5级D触发器
   pDFF dff4(ShReg[5], ShReg[4], Clock, Reset); // 第4级D触发器
   pDFF dff3(ShReg[4], ShReg[3], Clock, Reset); // 第3级D触发器
   pDFF dff2(ShReg[3], ShReg[2], Clock, Reset); // 第2级D触发器
   pDFF dff1(ShReg[2], ShReg[1], Clock, Reset); // 第1级D触发器
   pDFF dff0(ShReg[1], ShReg[0], Clock, Reset); // 第0级D触发器

   //===========================================================================
   // 奇偶校验运算
   // 对卷积结果的所有位进行异或运算，产生编码位
   //===========================================================================
   assign Yt[1] = wA[0] ^ wA[1] ^ wA[2] ^ wA[3] ^ wA[4] ^ wA[5] ^ wA[6] ^ wA[7] ^ wA[8];
   assign Yt[0] = wB[0] ^ wB[1] ^ wB[2] ^ wB[3] ^ wB[4] ^ wB[5] ^ wB[6] ^ wB[7] ^ wB[8];

   //===========================================================================
   // 输出同步
   // 将编码结果通过D触发器同步输出
   //===========================================================================
   pDFF dffy1(Yt[1], Y[1], Clock, Reset);     // 同步输出Y[1]
   pDFF dffy0(Yt[0], Y[0], Clock, Reset);     // 同步输出Y[0]

endmodule